`timescale 1ns / 1ps
module ins_decoder(
    input [31:0] ins,
    output reg [31:0] code
    );
    wire [5:0]   op;
    wire [5:0] func;
    assign op = ins[31:26];
    assign func = ins[5:0];

    always @(*)
    begin
        casez({op,func})
            //R-type
            12'b000000_100000:code <= 32'b00000000000000000000000000000001;//ADD   0
            12'b000000_100001:code <= 32'b00000000000000000000000000000010;//ADDU  1
            12'b000000_100010:code <= 32'b00000000000000000000000000000100;//SUB   2  
            12'b000000_100011:code <= 32'b00000000000000000000000000001000;//SUBU  3
            12'b000000_100100:code <= 32'b00000000000000000000000000010000;//AND   4
            12'b000000_100101:code <= 32'b00000000000000000000000000100000;//OR    5
            12'b000000_100110:code <= 32'b00000000000000000000000001000000;//XOR   6
            12'b000000_100111:code <= 32'b00000000000000000000000010000000;//NOR   7
            12'b000000_101010:code <= 32'b00000000000000000000000100000000;//SLT   8
            12'b000000_101011:code <= 32'b00000000000000000000001000000000;//SLTU  9
            12'b000000_000000:code <= 32'b00000000000000000000010000000000;//SLL   10
            12'b000000_000010:code <= 32'b00000000000000000000100000000000;//SRL   11
            12'b000000_000011:code <= 32'b00000000000000000001000000000000;//SRA   12
            12'b000000_000100:code <= 32'b00000000000000000010000000000000;//SLLV  13
            12'b000000_000110:code <= 32'b00000000000000000100000000000000;//SRLV  14
            12'b000000_000111:code <= 32'b00000000000000001000000000000000;//SRAV  15
            12'b000000_001000:code <= 32'b00000000000000010000000000000000;//JR    16
            //I-type
            12'b001000_??????:code <= 32'b00000000000000100000000000000000;//ADDI  17
            12'b001001_??????:code <= 32'b00000000000001000000000000000000;//ADDIU 18
            12'b001100_??????:code <= 32'b00000000000010000000000000000000;//ANDI  19
            12'b001101_??????:code <= 32'b00000000000100000000000000000000;//ORI   20
            12'b001110_??????:code <= 32'b00000000001000000000000000000000;//XORI  21
            12'b100011_??????:code <= 32'b00000000010000000000000000000000;//LW    22
            12'b101011_??????:code <= 32'b00000000100000000000000000000000;//SW    23
            12'b000100_??????:code <= 32'b00000001000000000000000000000000;//BEQ   24
            12'b000101_??????:code <= 32'b00000010000000000000000000000000;//BNE   25
            12'b001010_??????:code <= 32'b00000100000000000000000000000000;//SLTI  26
            12'b001011_??????:code <= 32'b00001000000000000000000000000000;//SLTIU 27
            12'b001111_??????:code <= 32'b00010000000000000000000000000000;//LUI   28
            12'b000010_??????:code <= 32'b00100000000000000000000000000000;//J     29
            12'b000011_??????:code <= 32'b01000000000000000000000000000000;//JAL   30
            default:          code <= 32'bx;
        endcase
    end 
endmodule
